LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY ProgramControler_Demo1 IS 
	PORT
	(
		CLOCK_50 :  IN  STD_LOGIC;
		KEY :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		SW :  IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX0 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX4 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX5 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX6 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX7 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		LEDG :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		LEDR :  OUT  STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END ProgramControler_Demo1;

ARCHITECTURE bdf_type OF ProgramControler_Demo1 IS 

COMPONENT programcontroller
	PORT(clk : IN STD_LOGIC;
		 programs_sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 state_in : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 temp_user_cook : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 temp_user_pre : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 time_user_cook : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 time_user_pre : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 out_desired_temp : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 out_desired_time : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT temperature_control
	PORT(clk : IN STD_LOGIC;
		 heat : IN STD_LOGIC;
		 cool : IN STD_LOGIC;
		 desired_temp_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 actual_temp_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT debounce
	PORT(clk : IN STD_LOGIC;
		 din : IN STD_LOGIC;
		 dout : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT timer
	PORT(enable : IN STD_LOGIC;
		 start : IN STD_LOGIC;
		 initial_val : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 done : OUT STD_LOGIC;
		 time_left : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bintobcd
	PORT(bin_input : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 bcd_output1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 bcd_output2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 bcd_output3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pulsegenerator
GENERIC (MAX : INTEGER
			);
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 pulse : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT button2
	PORT(CLK : IN STD_LOGIC;
		 PUSH_BUTTON_1 : IN STD_LOGIC;
		 PUSH_BUTTON_2 : IN STD_LOGIC;
		 out_temp : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT statemachine
	PORT(clk : IN STD_LOGIC;
		 timer_done : IN STD_LOGIC;
		 on_off : IN STD_LOGIC;
		 run : IN STD_LOGIC;
		 open_oven : IN STD_LOGIC;
		 enable7Seg : OUT STD_LOGIC;
		 starter_time : OUT STD_LOGIC;
		 food_in : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 state_out : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		 status : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pulsegenerator2
	PORT(clk : IN STD_LOGIC;
		 led_out : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT button
	PORT(CLK : IN STD_LOGIC;
		 PUSH_BUTTON_1 : IN STD_LOGIC;
		 PUSH_BUTTON_2 : IN STD_LOGIC;
		 out_temp : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT selectinput
	PORT(controle : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 entrada1 : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 entrada2 : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 saida : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ledblinker
	PORT(clk : IN STD_LOGIC;
		 led_out : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT enablecontrol
	PORT(enable : IN STD_LOGIC;
		 saida1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 saida2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT modeselector
	PORT(mode_sel : IN STD_LOGIC;
		 temp_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 time_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 temp_out_cook : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 temp_out_pre : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 time_out_cook : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 time_out_pre : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bin7segdecoder
	PORT(enable : IN STD_LOGIC;
		 binInput_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 binInput_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 binInput_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 decOut_0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 decOut_1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 decOut_2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT heatcool
	PORT(clk : IN STD_LOGIC;
		 state : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 heat : OUT STD_LOGIC;
		 cool : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT bin7segdecoder2
	PORT(enable : IN STD_LOGIC;
		 binInput_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 binInput_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 binInput_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 decOut_0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 decOut_1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(0 TO 8);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN 
SYNTHESIZED_WIRE_9 <= '1';
SYNTHESIZED_WIRE_12 <= '0';
SYNTHESIZED_WIRE_19 <= "111111111";



b2v_inst : programcontroller
PORT MAP(clk => CLOCK_50,
		 programs_sel => SW(5 DOWNTO 3),
		 state_in => SYNTHESIZED_WIRE_37,
		 temp_user_cook => SYNTHESIZED_WIRE_1,
		 temp_user_pre => SYNTHESIZED_WIRE_2,
		 time_user_cook => SYNTHESIZED_WIRE_3,
		 time_user_pre => SYNTHESIZED_WIRE_4,
		 out_desired_temp => SYNTHESIZED_WIRE_7,
		 out_desired_time => SYNTHESIZED_WIRE_10);


b2v_inst1 : temperature_control
PORT MAP(clk => CLOCK_50,
		 heat => SYNTHESIZED_WIRE_5,
		 cool => SYNTHESIZED_WIRE_6,
		 desired_temp_in => SYNTHESIZED_WIRE_7,
		 actual_temp_out => SYNTHESIZED_WIRE_27);


b2v_inst10 : debounce
PORT MAP(clk => CLOCK_50,
		 din => SW(0),
		 dout => SYNTHESIZED_WIRE_14);


b2v_inst11 : timer
PORT MAP(enable => SYNTHESIZED_WIRE_8,
		 start => SYNTHESIZED_WIRE_9,
		 initial_val => SYNTHESIZED_WIRE_10,
		 done => SYNTHESIZED_WIRE_13,
		 time_left => SYNTHESIZED_WIRE_11);


b2v_inst13 : bintobcd
PORT MAP(bin_input => SYNTHESIZED_WIRE_11,
		 bcd_output1 => SYNTHESIZED_WIRE_34,
		 bcd_output2 => SYNTHESIZED_WIRE_35,
		 bcd_output3 => SYNTHESIZED_WIRE_36);


b2v_inst14 : pulsegenerator
GENERIC MAP(MAX => 50000000
			)
PORT MAP(clk => CLOCK_50,
		 reset => SYNTHESIZED_WIRE_12,
		 pulse => SYNTHESIZED_WIRE_8);



b2v_inst16 : debounce
PORT MAP(clk => CLOCK_50,
		 din => SW(1),
		 dout => SYNTHESIZED_WIRE_15);


b2v_inst17 : debounce
PORT MAP(clk => CLOCK_50,
		 din => SW(2),
		 dout => SYNTHESIZED_WIRE_16);


b2v_inst2 : button2
PORT MAP(CLK => CLOCK_50,
		 PUSH_BUTTON_1 => KEY(2),
		 PUSH_BUTTON_2 => KEY(3),
		 out_temp => SYNTHESIZED_WIRE_25);


b2v_inst22 : statemachine
PORT MAP(clk => CLOCK_50,
		 timer_done => SYNTHESIZED_WIRE_13,
		 on_off => SYNTHESIZED_WIRE_14,
		 run => SYNTHESIZED_WIRE_15,
		 open_oven => SYNTHESIZED_WIRE_16,
		 enable7Seg => SYNTHESIZED_WIRE_38,
		 food_in => SYNTHESIZED_WIRE_17,
		 state_out => SYNTHESIZED_WIRE_37,
		 status => SYNTHESIZED_WIRE_23);


LEDG <= SYNTHESIZED_WIRE_17 AND SYNTHESIZED_WIRE_18;


b2v_inst28 : pulsegenerator2
PORT MAP(clk => CLOCK_50,
		 led_out => SYNTHESIZED_WIRE_18);


b2v_inst3 : button
PORT MAP(CLK => CLOCK_50,
		 PUSH_BUTTON_1 => KEY(0),
		 PUSH_BUTTON_2 => KEY(1),
		 out_temp => SYNTHESIZED_WIRE_26);


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20;


b2v_inst32 : selectinput
PORT MAP(controle => SYNTHESIZED_WIRE_37,
		 entrada1 => SYNTHESIZED_WIRE_22,
		 entrada2 => SYNTHESIZED_WIRE_23,
		 saida => LEDR);


b2v_inst33 : ledblinker
PORT MAP(clk => CLOCK_50,
		 led_out => SYNTHESIZED_WIRE_20);



b2v_inst37 : enablecontrol
PORT MAP(enable => SYNTHESIZED_WIRE_38,
		 saida1 => HEX4,
		 saida2 => HEX5);


b2v_inst4 : modeselector
PORT MAP(mode_sel => SW(6),
		 temp_in => SYNTHESIZED_WIRE_25,
		 time_in => SYNTHESIZED_WIRE_26,
		 temp_out_cook => SYNTHESIZED_WIRE_1,
		 temp_out_pre => SYNTHESIZED_WIRE_2,
		 time_out_cook => SYNTHESIZED_WIRE_3,
		 time_out_pre => SYNTHESIZED_WIRE_4);


b2v_inst5 : bintobcd
PORT MAP(bin_input => SYNTHESIZED_WIRE_27,
		 bcd_output1 => SYNTHESIZED_WIRE_29,
		 bcd_output2 => SYNTHESIZED_WIRE_30,
		 bcd_output3 => SYNTHESIZED_WIRE_31);


b2v_inst6 : bin7segdecoder
PORT MAP(enable => SYNTHESIZED_WIRE_38,
		 binInput_0 => SYNTHESIZED_WIRE_29,
		 binInput_1 => SYNTHESIZED_WIRE_30,
		 binInput_2 => SYNTHESIZED_WIRE_31,
		 decOut_0 => HEX0,
		 decOut_1 => HEX1,
		 decOut_2 => HEX2);


b2v_inst7 : heatcool
PORT MAP(clk => CLOCK_50,
		 state => SYNTHESIZED_WIRE_37,
		 heat => SYNTHESIZED_WIRE_5,
		 cool => SYNTHESIZED_WIRE_6);


b2v_inst8 : bin7segdecoder2
PORT MAP(enable => SYNTHESIZED_WIRE_38,
		 binInput_0 => SYNTHESIZED_WIRE_34,
		 binInput_1 => SYNTHESIZED_WIRE_35,
		 binInput_2 => SYNTHESIZED_WIRE_36,
		 decOut_0 => HEX6,
		 decOut_1 => HEX7);



END bdf_type;